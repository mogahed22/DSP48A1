module DSP48A1(
    AIN,BIN,CIN,DIN,OPMODEIN,PCIN,CARRYININ,BCIN,PCLK,PCE,PRST,
    BCOUT,M,CARRYOUTOUT,CARRYOUTOUTOFF,P,PCOUT,XIN0,ZIN0
    ); 

//parameters 
parameter SYNCD = 1'b0;
parameter ASYNCD = 1'b1;
parameter RSTTYPED = SYNCD ;
parameter A0REGD = 0 ;
parameter A1REGD = 1;
parameter B0REGD = 0;
parameter B1REGD = 1;
parameter DIRECTIOND = "DIRECT";
parameter CREGD = 1;
parameter DREGD = 1;
parameter PREGD = 1;
parameter CARRYOUTREGD = 1;
parameter CARRYINREGD = 1;
parameter OPMODEREGD = 1;
parameter MREGD = 1;

parameter CARRYINSEL = "OPMODE5";

//inputs decleration
input [17:0] AIN,BIN,DIN,BCIN;
input [47:0] CIN,PCIN;
input [7:0] OPMODEIN;
input CARRYININ,PCLK,PCE,PRST;
input [47:0] XIN0 = 0; 
input[47:0] ZIN0 =0;

//outputs decleration
output [47:0] P,PCOUT;
output [35:0] M;
output [17:0] BCOUT;
output CARRYOUTOUT,CARRYOUTOUTOFF;

//wires decleration
wire [17:0] DO , B0O , PRASO , MUXYO , B1O , A0O , A1O ;
wire [47:0] CO,MULTIPLYERO , MREGO ,  XOUT , DAB , PX , PZ , ZOUT ;
wire [48:0] PTSAO;
wire [7:0] OPMODEO;
wire CARRYCASCADE , CARRYINOUT;


//Moduls instantiations 
OPMODEREG #(.SYNC(SYNCD),.ASYNC(ASYNCD),.RSTTYPE(RSTTYPED),.OPMODEREG(OPMODEREGD))opmodereg (
    .OPMODE(OPMODEIN),.OPMODE_mux(OPMODEO),.CLK(PCLK),.CEOPMODE(PCE),.RSTOPMODE(PRST));

DREG #(.SYNC(SYNCD),.ASYNC(ASYNCD),.RSTTYPE(RSTTYPED),.DREG(DREGD)) dreg(
    .D(DIN),.Dmux(DO),.CLK(PCLK),.RSTD(PRST),.CED(PCE));

B0REG #(.SYNC(SYNCD),.ASYNC(ASYNCD),.RSTTYPE(RSTTYPED),.B0REG(B0REGD)) b0reg(
    .BINPUT(BIN),.BCASCADED(BCIN),.B_mux0(B0O),.CLK(PCLK),.RSTB(PRST),.CEB(PCE));

B1REG #(.SYNC(SYNCD),.ASYNC(ASYNCD),.RSTTYPE(RSTTYPED),.B1REG(B1REGD)) b1reg(
    .B1(MUXYO),.B_mux1(B1O),.CLK(PCLK),.RSTB(PRST),.CEB(PCE));

A0REG #(.SYNC(SYNCD),.ASYNC(ASYNCD),.RSTTYPE(RSTTYPED),.A0REG(A0REGD)) a0reg (
    .A0(AIN),.A_mux0(A0O),.CLK(PCLK),.RSTA(PRST),.CEA(PCE));

A1REG #(.SYNC(SYNCD),.ASYNC(ASYNCD),.RSTTYPE(RSTTYPED),.A1REG(A1REGD)) a1reg(
    .A1(A0O),.A_mux1(A1O),.CLK(PCLK),.RSTA(PRST),.CEA(PCE));

MREG #(.SYNC(SYNCD),.ASYNC(ASYNCD),.RSTTYPE(RSTTYPED),.MREG(MREGD)) mreg (
    .M(MULTIPLYERO),.M_mux(MREGO),.CLK(PCLK),.RSTM(PRST),.CEM(PCE));

CREG #(.SYNC(SYNCD),.ASYNC(ASYNCD),.RSTTYPE(RSTTYPED),.CREG(CREGD)) creg (
    .C(CIN),.Cmux(CO),.CLK(PCLK),.RSTC(PRST),.CEC(PCE));

CARRYINREG #(.SYNC(SYNCD),.ASYNC(ASYNCD),.RSTTYPE(RSTTYPED),.CARRYINREG(CARRYINREGD)) carryinreg(
    .CARRYIN(CARRYCASCADE),.CARRYIN_mux(CARRYINOUT),.CLK(PCLK),.RSTCARRYIN(PRST),.CECARRYIN(PCE));

CARRYOUTREG #(.SYNC(SYNCD),.ASYNC(ASYNCD),.RSTTYPE(RSTTYPED),.CARRYOUTREG(CARRYOUTREGD)) carryoutreg(
    .CARRYOUT(PTSAO[48]),.CARRYOUT_mux(CARRYOUTOUT),.CLK(PCLK),.RSTCARRYIN(PRST),.CECARRYIN(PCE));

PREG #(.SYNC(SYNCD),.ASYNC(ASYNCD),.RSTTYPE(RSTTYPED),.PREG(PREGD)) preg(
    .P(PTSAO[47:0]),.P_mux(P),.CLK(PCLK),.RSTP(PRST),.CEP(PCE));


assign PX = P;
assign PZ = P;
//assign XIN0 =48'b0;
//assign ZIN0 =48'b0;
assign DAB = {DO[11:0],A1O[17:0],B1O[17:0]};
assign PRASO = (OPMODEO[6]) ? B0O+DO : DO-B0O;
assign MUXYO = (OPMODEO[4]) ? PRASO : B0O;
assign MULTIPLYERO = B1O * A1O ;
assign M = MREGO [35:0];
assign BCOUT = B1O;
assign XOUT= (OPMODEO[1:0]==0)? 48'b0 : (OPMODEO[1:0] == 1)? MREGO :(OPMODEO[1:0] == 2)? PX :(OPMODEO[1:0]==3)? DAB : 48'b0;
assign ZOUT = (OPMODEO[3:2]==0)? 48'b0 :(OPMODEO[3:2]==1)? PCIN :(OPMODEO[3:2]==2)? PZ:(OPMODEO==3)? CO :48'b0;
assign CARRYCASCADE = (CARRYINSEL=="OPMODE5")? OPMODEO[5] :(CARRYINSEL=="CARRYIN")?CARRYININ : 1'b0;
assign PTSAO[47:0] = (OPMODEO[7]==0)? XOUT + ZOUT :(OPMODEO[7]==1)? ZOUT-(XOUT+CARRYINOUT) :48'b0;
assign CARRYOUTOUTOFF = CARRYOUTOUT;
assign PCOUT = P;


endmodule